module ProgramCounter(AddressMux, address);
//initialize size of address 
parameter SIZE = 5;

//initialize port
input[SIZE-1:0] AddressMux;
output reg[SIZE-1:0] address;



endmodule
